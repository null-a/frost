`default_nettype none

module top (input clk);
endmodule // top
