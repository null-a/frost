`default_nettype none

module fpga_tb();
endmodule // fpga_tb
